//0416221 劉川楓, 0416251 梁幸儀
//Subject:     CO project 2 - Sign extend
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Sign_Extend(
    data_i,
	isORI_i,
    data_o
    );
               
//I/O ports
input   [16-1:0] data_i;
input   isORI_i;
output  [32-1:0] data_o;

//Internal Signals
reg     [32-1:0] data_o;



//Sign extended
always@(*) begin
	data_o[15:0]<=data_i;
	if(data_i[15] == 0 || isORI_i)
		data_o[31:16]<=16'b0000000000000000;
	else
		data_o[31:16]<=16'b1111111111111111;
end
endmodule      
     